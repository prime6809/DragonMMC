`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:			Ramoth 
// Engineer: 		Phill Harvey-Smith.
// 
// Create Date:    	15:57:34 06/29/2011 
// Design Name: 	DragonMMC
// Module Name:    	Main 
//
// **NOTE** if source looks oddly formatted in ISE, set editor tab width to 4!
//
//////////////////////////////////////////////////////////////////////////////////
//
// Dragon 		Dir		Function
// address	
//
// $FF50		R		AVR Result
// $FF50		 W		AVR command
// $FF51		 W		AVR 'latch' reg for single byte params.
// $FF52		R		AVR Read data register
// $FF53		 W		AVR Write data register
// $FF54		R		AVR Status, busy etc, handshake bits
// $FF55		 W		PIA redirect if b0 written 1.
// $FF56		RW		RAM / ROM control register
// $FF57 unused?
// $FF58		R		Sam bits MSB
// $FF59		R		Sam bits LSB
// $FF5A		RW		RAM bank for RAM reads
// $FF5B		RW		RAM bank for RAM writes
// $FF5C unused
// $FF5D unused
// $FF5E unused
// $FF5F unused
//
// **Note** throughout the module I use positive logic, and then invert before 
// driving the output if needed. I do this as then I know that I can do 
// if (signal) and it has an unambiguous meaning. 
//

module DragonMMC(
	// 6809 side
    input [15:0] Addr,		// Dragon address bus
    inout [7:0] Data,		// Daragon data bus
    input E,				// E clock
	input Q,				// Q clock
    input RW,				// Read/Write
    input CSEL,				// Cart rom select 
    input P2,				// P2/SCS acrive from $ff40-$ff5f
    input Reset,			// System reset
	output DSD,				// Device select disable
    output CART,			// Cart FIRQ
    output NMI,				// Non maskable interupt
    output HALT,			// Halt CPU
    
	// AVR side 
    inout [7:0] AData,		// AVR data bus
    input [1:0] AAddr,		// AVR data bus
    input nARD,				// AVR read strobe
    input nAWR,				// AVR write strobe
    input AVRBusy,			// AVR busy when 1
	output AInt,			// Interupt to AVR
	
	// Memory control
    output nRD,				// Read strobe
    output nWR,				// Write strobe
    output nROMCS,			// ROM chip select
    output nRAMCS,			// RAM chip select
	output reg ROMA14,		// A14 pin for rom, used to select between Dragon(0) & CoCo(1) versions of ROM
	output [18:15] RAMA,	// RAM upper address lines.
	
	// Snapshot button
	input	ANMI,			// AVR NMI generated by Snapshot button 
	
	// Force Cold reset button
	input	nFCReset,		//  Button on board, when pressed along with reset, forces back to rom mode.
	
	// Spare pins currently unassigned.
	inout [8:0] SP,
	inout Pin2,
	inout Pin7,
	inout Pin46,
	inout Pin80,
	inout Pin85,
		
	// I/O Port, currently unused.
    inout [7:0] FData		// FTDI data bus
    );

	
	// Memory Mapping bits

	reg		RamEnable;		// Should RAM be ebnabled in the $8000-$FEFF area ?
	reg		PIAReg;			// Should we replace PIA data at $FF20 ?
	reg		RAMVec;			// Should we read interrupt vectors from ROM or RAM
	
	// 6809 and AVR output data registers.
	
	reg [7:0] 	DragonToAVR;	// Data going from Dragon -> AVR
	reg [7:0] 	AVRToDragon;	// Data going from AVR -> Dragon
	reg [3:0]	AddrLatch;		// Latch of written address. (This could be reduced to 2 bits - PHS 2017-04-04).
	reg 		DragonRW;		// Did the dragon read or write ?
	reg			RamWP;			// Ram Write protect
	reg			RomWE;			// EEPROM write enable.
	reg			FIRQEn;			// FIRQ routing enable

	reg	[3:0]	RamRPtr = 4'b0;		// RAM Read bank pointer
	reg	[3:0]	RamWPtr = 4'b0;		// RAM Write bank pointer

	// Handshake bits
	reg			DragonW_AVRR;	// Set by Dragon write, cleared by AVR read.
	reg			AVRW_DragonR;	// Set by AVR write, cleared by Dragon read.
	reg			NMIEn;			// Set if NMI from AVR enabled.
	reg			IntRAMWP;		// Interrupt area RAM write protect

	reg	[15:0]	SAMBits ;		// 1 bit x 16 bit array.....
	
	// Previously this was a seperate latch.
	assign	MapMode		= SAMBits[15];

	reg		MotorON;			// Captured motor control bit
	
// If NMI is enabled, it will follow the ANMI line, otherwise let it float high 

	assign NMI			= NMIEn ? ANMI : 1'bz;

// Not used currently so set to zero for compatibility.....
//	assign RAMA[18:15]	= 4'b0000;

	// Generate OE and WE signals, only do this if Reset is high ! 
	assign RD			= E & RW & Reset;
	assign WR			= E & ~RW & Reset;
	assign nRD			= ~RD;
	assign nWR			= ~WR; 


// Cold reset signal high only if reset low *AND* ColdReset button pressed. 
// This allows us to get back to the onboard ROMs without having to powercycle.
// if we have loaded a Cartridge image into the $C000-$FEFF area.
	assign ColdReset	= (Reset | nFCReset) == 1'b0;

//
// Address decoding and ROM/RAM banking control.
// 	
	
	// Memory control register as follows :
	// 
	// Bit		Function
	// 0		When 1 enable the RAM between $8000 and $FEFF for both reads and writes, disables internal and cart ROMS.
	// 1		When 1 write protect the rom once enabled.
	// 2		When 1 enable routing of the Q signal to the FIRQ line, to auto-start the cartridge (normally an image in RAM).
	// 3		When 1 enable writes to the EEPROM/Flash, so that it can be updated (if jumper set to WE position).
	// 4		Routed to line A14 of the EEPROM/Flash, to select either Dragon (0) or CoCo (1) version of the firmware.
	// 5		When 1 Read interrupt vectors from RAM, otherwise ROM as normal
	// 6		When 1 pressing Snap button on AVR will generate an NMI on 6809.
	// 7		When 1 Interrupt area RAM is write protected.
	//
	assign RamCTRL		= (Addr==16'hFF56);
	assign RamCTRLRD	= RamCTRL & RD;
	assign RamCTRLWR	= RamCTRL & WR;
	
	always @(negedge RamCTRLWR or posedge ColdReset)
	begin
		if (ColdReset) 
		begin
			RamEnable	<= 1'b0;
			RamWP		<= 1'b0;
			FIRQEn		<= 1'b0;
			RomWE		<= 1'b0;
			ROMA14		<= 1'b0;
			RAMVec		<= 1'b1;
			NMIEn		<= 1'b1;
			IntRAMWP	<= 1'b1;
		end
		else
		begin
			RamEnable	<= Data[0];
			RamWP		<= Data[1];
			FIRQEn		<= Data[2];
			RomWE		<= Data[3];
			ROMA14		<= Data[4];
			RAMVec		<= Data[5];
			NMIEn		<= Data[6];
			IntRAMWP	<= Data[7];
		end
	end
	
	// Ram Read and write bank registers.
	// Write / Reset control.
	assign RamRPtrEn	= (Addr==16'hFF5A);
	assign RamRPtrRE	= RamRPtrEn & RD;
	assign RamRPtrWE	= RamRPtrEn & WR;
	
	assign RamWPtrEn	= (Addr==16'hFF5B);
	assign RamWPtrRE	= RamWPtrEn & RD;
	assign RamWPtrWE	= RamWPtrEn & WR;
	
	always @(negedge RamRPtrWE or negedge Reset)
	begin
		if (!Reset)
			RamRPtr	<= 4'b0000;
		else
			RamRPtr	<= Data[3:0];
	end
	
	always @(negedge RamWPtrWE or negedge Reset)
	begin
		if (!Reset)
			RamWPtr	<= 4'b0000;
		else
			RamWPtr	<= Data[3:0];
	end
	
	// PIA replace register, write only!
	assign PIAReplace	= (Addr==16'hFF55) & WR;
	
	// Bottom bit written latched directly into PIA control latch
	always @(negedge PIAReplace or negedge Reset)
	begin
		if (!Reset)
			PIAReg 	<= 1'b0;
		else
			PIAReg	<= Data[0];
	end
	
	
	// CART/FIRQ redirect Q to CART if enabled. This allows loaded cartridge
	// images to auto-start like a normal game cartridge.
	assign CART		= FIRQEn ? Q : 1'bz;
	
	// Address ranages
	assign RangeRAM		= ((Addr>=16'h8000) && (Addr<=16'hFEFF));
	assign RangeROM		= ((Addr>=16'hC000) && (Addr<=16'hFEFF));
	assign RangePIA		= (Addr==16'hFF20);
	assign RangeMotor	= (Addr==16'hFF21);
	
	// 14 bytes of vectors + 2 bytes 'reserved', was previously FFE0 and above, but this
	// clashes with the DragonPlus board which uses FFE0-FFE2.
	assign RangeInt		= ((Addr>=16'hFFF0) && (Addr<=16'hFFFF));		
	
	assign RomRead		= RangeROM & RD & ~RamEnable & ~MapMode;
	assign RomWrite		= RangeROM & WR & RomWE & ~RamEnable & ~MapMode;
	
	assign RamRead		= RangeRAM & RD & RamEnable & ~MapMode;
	assign RamWrite		= RangeRAM & WR & ~RomWE & ~RamWP & ~MapMode;
		
	assign IntRead		= RangeInt & RD & RAMVec;
	assign IntWrite		= RangeInt & WR & ~RomWE & ~IntRAMWP;
	
	// Enable ROM if we are in map mode 0 and RamEnable is false.
	assign ROMCS		= RomRead | RomWrite;
	assign nROMCS		= ~ROMCS;

	// Enable ram either when writing to the RAM range or when reading from the range with 
	// RamEnable set, this way writes always go to the RAM.
	// 2016-04-05, ram disabled if writing and RomWE is set, for update of ROM.
	// Do not enable the RAM in MapMode 1 as onboard RAM enabled then.
	// Enable top 16 bytes of RAM if writing to vectors, or reading them from RAM (default is from ROM).
	assign RAMCS		= RamRead | RamWrite | IntRead | IntWrite;
	assign nRAMCS		= ~RAMCS;
	assign RAMA[18:15]	= RangeInt ? 4'b0000 : 
						  RamWrite ? RamWPtr[3:0] : RamRPtr[3:0];

	// Enable signal if we are replacing PIA reg at $FF20 for tape emulation.
	assign PIACS		= RangePIA & PIAReg & RD;
	assign nPIACS		= ~PIACS;
//
// AVR<-->Dragon data exchange
//
	assign DragonIO		= ((Addr>=16'hff50) && (Addr<=16'hff53));
	assign DragonIORD	= DragonIO & RD;
	assign DragonIOWR	= DragonIO & WR;
	
	assign AVRStatus	= (Addr == 16'hff54);		// AVR status at $FF54
	assign AVRStatusRD	= AVRStatus & RD;

//
// Capture writes to the 16 SAM 'registers'.
//
// The SAM has 16 configuration bits which are cleared by writing to an even address
// and written by writing to an odd address. These are mapped in between $FFC0 and 
// $FFDF. The reason for this is that the SAM does not have a connection to the data
// bus due to a lack of package pins.
// We can capture this information by triggering a latch of the bottom address bit 
// when a write is made to this range and using address bits 4..1 (effectively) 
// shifted left one bit as an index to the array of bits.
// 
	assign SAMBitsAddr	= ((Addr>=16'hFFC0) && (Addr<=16'hFFDF));
	assign SAMBitsWR	= SAMBitsAddr & WR;
	
	wire [3:0] SAMReg;
	assign SAMReg[3:0]	= Addr[4:1];
	
	always @(posedge SAMBitsWR or negedge Reset)
	begin
	  if (!Reset)
	  begin
        SAMBits[15:0] <= 16'h0000;
	  end
	  else
	  begin
        SAMBits[SAMReg[3:0]] <= Addr[0];
	  end
	end

//
// Output SAM bits in 2 consecutive 6809 memory locations, that way we can do a 
// 16 bit read to get them all in one go.
//	
	assign SAMBitsH		= (Addr==16'hFF58);
	assign SAMBitsL		= (Addr==16'hFF59);
	
	assign SAMBitsRD	= (SAMBitsL | SAMBitsH) & RD;

	wire [7:0]	SAMData;
	assign SAMData		= SAMBitsL ? SAMBits[7:0] : SAMBits[15:8];

	assign AddrLatchEN	= DragonIOWR; 
	assign AInt			= DragonIORD | DragonIOWR;

	// Capture the bottom 4 address lines on a write by the Dragon to our IO registers
	// or to one ofg the SAM registers
	// 2017-04-04, PHS, since the AVR registers only span 4 locations and the AVR is 
	// no longer handling SAM bit writes, this should be able to be reduced to 2 bits.
	always @(posedge AddrLatchEN or negedge Reset)
	begin
	  if(!Reset)
	  begin
	    AddrLatch[3:0] <= 4'b0000;
	  end
	  else
	  begin
	    AddrLatch[3:0] <= Addr[3:0];
	  end
	end

	// Latch read or write
	always @(posedge AInt)
	begin
	  DragonRW <= RW;
	end

	// When the AVR reads give it the Dragon data / latched address
	wire [7:0]	AVRDataOut;
	assign 	AVRDataOut[7:0]	= AAddr[0] ? { MotorON, DragonRW,2'b0,AddrLatch[3:0] } : DragonToAVR[7:0];
	assign	AData			= nARD ? 8'bz : AVRDataOut;
	
	// When the Dragon reads give it the AVR data / status
	// Note both reading the AVR data reg & the PIA override give the AVRToDragon reg.
	wire [7:0] 	DragonDataOut;
	assign 	DragonDataOut[7:0]		= 
									  RamRPtrRE ? {4'b0,RamRPtr } :
									  RamWPtrRE ? {4'b0,RamWPtr } :
									  SAMBitsRD ? SAMData :
									  AVRStatus ? {5'b0,AVRW_DragonR,DragonW_AVRR,AVRBusy} : 
									  RamCTRLRD	? {IntRAMWP,NMIEn,RAMVec,ROMA14, RomWE, FIRQEn, RamWP, RamEnable} :
											AVRToDragon;
	
	assign 	Data					= (DragonIORD | AVRStatusRD | RamCTRLRD | SAMBitsRD | PIACS | RamRPtrRE | RamWPtrRE) ? DragonDataOut : 8'bz;
//	assign 	Data					= (DragonIORD | AVRStatusRD | RamCTRLRD | SAMBitsRD | PIACS ) ? DragonDataOut : 8'bz;

	assign 	FData					= {5'b0,AVRW_DragonR,DragonW_AVRR,AVRBusy};
	
	// Latch Dragon to AVR reg on Dragon write
	always @(negedge DragonIOWR)
	begin
	  DragonToAVR <= Data;
	end
	
	// Latch AVR to Dragon on AVR write
	always @(negedge nAWR)
	begin
	  AVRToDragon <= AData;
	end
	
	// Handshake lines.
	// DragonW_AVRR set by a write from the Dragon, cleared by a read by the AVR.
	// Cleared on reset.
	always @(negedge Reset or posedge DragonIOWR or negedge nARD)
	begin
		if(!Reset)
			DragonW_AVRR <= 1'b0;
		else if(DragonIOWR)
			DragonW_AVRR <=  1'b1;
		else
			DragonW_AVRR <= 1'b0;
	end

	// AVRW_DragonR set by a write from the AVR, cleared by a read by the Dragon.
	// Cleared on reset.
	always @(negedge Reset or posedge DragonIORD or negedge nAWR)
	begin
		if(!Reset)
			AVRW_DragonR <= 1'b0;
		else if(DragonIORD)
			AVRW_DragonR <=  1'b0;
		else
			AVRW_DragonR <= 1'b1;
	end
	
	// 
	// Capture bit 3 of writes to PIA1 control register A, as this controls the
	// cassette motor.
	//
	
	assign MotorWR	= RangeMotor & WR;
	
	always @(negedge Reset or negedge MotorWR)
	begin
	  if(!Reset)
	    MotorON <= 1'b0;
	  else
	    MotorON <= Data[3];
	end
	
	
	// Disable internal device selection only when our ram or I/O is enabled
	// or we are replacing PIA reg.
	assign DSD			= (RAMCS | PIACS | DragonIO | AVRStatus | PIAReplace | RamCTRL | SAMBitsH | SAMBitsL | RamRPtrEn | RamWPtrEn) ? 1'b0 : 1'bz;
	
	assign HALT = 1'bz;
endmodule
